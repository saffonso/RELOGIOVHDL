library verilog;
use verilog.vl_types.all;
entity Relogio_vlg_vec_tst is
end Relogio_vlg_vec_tst;
